library verilog;
use verilog.vl_types.all;
entity monitor_tb is
end monitor_tb;
