module div_3(
    input clk,
    input [7:0] in,
    output reg [7:0] out
);


endmodule
