module top(
    input CLOCK_50,
    output [7:0] LEDG,
    output [9:5] LEDR,
    output [6:0] HEX3,
    output [6:0] HEX2,
    output [6:0] HEX1,
    output [6:0] HEX0,
    output [11:0] DRAM_ADDR,
    output DRAM_BA_1,
    output DRAM_BA_0,
    output DRAM_CAS_N,
    output DRAM_RAS_N,
    output DRAM_CLK,
    output DRAM_CKE,
    output DRAM_CS_N,
    output DRAM_WE_N,
    output DRAM_UDQM,
    output DRAM_LDQM,
    inout [15:0] DRAM_DQ
);

    wire toggle_clock;
    nios_system u0 (
        .green_leds_external_connection_export (LEDG), // green_leds_external_connection.export
        .hex3_external_connection_export       (HEX3),       //       hex3_external_connection.export
        .hex2_external_connection_export       (HEX2),       //       hex2_external_connection.export
        .hex1_external_connection_export       (HEX1),       //       hex1_external_connection.export
        .hex0_external_connection_export       (HEX0),       //       hex0_external_connection.export
        .altpll_0_inclk_interface_clk          (CLOCK_50),          //       altpll_0_inclk_interface.clk
        .altpll_0_c2_clk                       (toggle_clock),                       //                    altpll_0_c2.clk
        .clock_bridge_0_out_clk_1_clk          (DRAM_CLK),          //       clock_bridge_0_out_clk_1.clk
        .sdram_0_wire_addr                     (DRAM_ADDR),                     //                   sdram_0_wire.addr
        .sdram_0_wire_ba                       ({DRAM_BA_1, DRAM_BA_0}),                       //                               .ba
        .sdram_0_wire_cas_n                    (DRAM_CAS_N),                    //                               .cas_n
        .sdram_0_wire_cke                      (DRAM_CKE),                      //                               .cke
        .sdram_0_wire_cs_n                     (DRAM_CS_N),                     //                               .cs_n
        .sdram_0_wire_dq                       (DRAM_DQ),                       //                               .dq
        .sdram_0_wire_dqm                      ({DRAM_UDQM, DRAM_LDQM}),                      //                               .dqm
        .sdram_0_wire_ras_n                    (DRAM_RAS_N),                    //                               .ras_n
        .sdram_0_wire_we_n                     (DRAM_WE_N)                      //                               .we_n
    );

    toggle t(toggle_clock, LEDR);

endmodule

module toggle(
    input clk,
    output [9:5] counter_out
);

    reg [31:0] counter_data;

    always @(posedge clk)
        counter_data <= counter_data + 1;

    assign counter_out[9] = counter_data[21];
    assign counter_out[5] = counter_data[21];
    assign counter_out[8] = counter_data[26];
    assign counter_out[6] = counter_data[26];
    assign counter_out[7] = counter_data[27];

endmodule
